//=============================================================================
// Project       : AXI VIP
//=============================================================================
// Filename      : axi_timescale.sv
// Author        : VLSI GROUP
// Company       : NO
// Date          : 03-Jan-2022
//=============================================================================
// Description   : 
//
//
//
//=============================================================================
`ifndef GUARD_AXI_TIMESCALE__SV
`define GUARD_AXI_TIMESCALE__SV

timeunit 1ps;
timeprecision 1ps;

`endif


