//=============================================================================
// Project       : AXI VIP
//=============================================================================
// Filename      : axi_if.sv
// Author        : VLSI GROUP
// Company       : NO
// Date          : 03-Jan-2022
//=============================================================================
// Description   : 
//
//
//
//=============================================================================
`ifndef GUARD_AXI_IF__SV
`define GUARD_AXI_IF__SV

interface axi_if();

  logic  aclk;   
  logic  aresetn;

endinterface

`endif


