package vt_axi_pkg;
  struct {
    logic 
  } awaddr_s

endpackage