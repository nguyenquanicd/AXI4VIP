//=============================================================================
// Project       : AXI VIP
//=============================================================================
// Filename      : axi_test_pkg.sv
// Author        : VLSI GROUP
// Company       : NO
// Date          : 03-Jan-2022
//=============================================================================
// Description   : 
//
//
//
//=============================================================================
`ifndef GUARD_AXI_TEST_PACKAGE__SV
`define GUARD_AXI_TEST_PACKAGE__SV

package axi_test_pkg;
  import uvm_pkg::*;

  import axi_pkg::*;
  import axi_sequence_pkg::*;
  import axi_environment_pkg::*;

  `include "axi_base_test.sv";

endpackage: axi_test_pkg

`endif


